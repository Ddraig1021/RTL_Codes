LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CLOCK_DIVIDER IS
	PORT
	(
		SYS_CLK : IN STD_LOGIC;
		CLK_OUT : OUT STD_LOGIC 
	);
END CLOCK_DIVIDER;

ARCHITECTURE RTL OF CLOCK_DIVIDER IS
	SIGNAL COUNTER : INTEGER := 0 TO 10 := 0;
	SIGNAL TOGGLE : STD_LOGIC := '0';
BEGIN  
PROCESS(SYS_CLK)
BEGIN
	IF RISING_EDGE(SYS_CLK) THEN 
		IF COUNTER = 9 THEN
			COUNTER <= 0;
			TOGGLE <= NOT TOGGLE;
		ELSE
			COUNTER <= COUNTER + 1;
		END IF;
	END IF;
END PROCESS;

CLK_OUT <= TOGGLE;

END RTL;